**SRAM
Vd 3 0 dc 5v
Vq 1 0 dc 0v
Vqb 2 0 dc 5v
Vw 4 0 pulse(5 0 0 0 0 50ms 100ms)
C1 5 0 0.1p
C2 6 0 0.1p
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
m1 1 2 3 3 pmod w=100u l=10u
m2 1 2 0 0 nmod w=100u l=10u
m3 2 1 3 3 pmod w=100u l=10u
m4 2 1 0 0 nmod w=100u l=10u
m5 1 4 5 0 nmod w=100u l=10u
m6 2 4 6 0 nmod w=100u l=10u
.tran 0.01ms 200ms
.control
run
plot V(4)
plot V(5)
plot V(6)
.endc
.end
