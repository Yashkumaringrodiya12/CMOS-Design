** Full adder using cmos technology
.subckt inverter 1 2 3
mp 2 1 3 3 pmod w=100u l=10u
mn 2 1 0 0 nmod w=100u l=10u
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
.ends
Vd 1 0 dc 5v
Va 11 0 pulse(0 5 0 0 0 10m 20m)
Vb 12 0 pulse(0 5 0 0 0 20m 40m)
Vci 13 0 pulse(0 5 0 0 0 40m 80m)
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
m1 14 12 0 0 nmod w=100u l=10u
m2 15 11 14 0 nmod w=100u l=10u
m3 16 12 0 0 nmod w=100u l=10u
m4 16 11 0 0 nmod w=100u l=10u
m5 15 13 16 0 nmod w=100u l=10u
m6 15 11 17 1 pmod w=100u l=10u
m7 15 12 17 1 pmod w=100u l=10u
m8 17 13 1 1 pmod w=100u l=10u
m9 18 11 1 1 pmod w=100u l=10u
m10 17 12 18 1 pmod w=100u l=10u
m11 18 11 0 0 nmod w=100u l=10u
m12 18 12 0 0 nmod w=100u l=10u
m13 18 13 0 0 nmod w=100u l=10u
m14 19 13 0 0 nmod w=100u l=10u
m15 20 12 19 0 nmod w=100u l=10u
m16 21 11 20 0 nmod w=100u l=10u
m17 21 15 18 0 nmod w=100u l=10u
m18 21 11 22 1 pmod w=100u l=10u
m19 21 12 22 1 pmod w=100u l=10u
m20 21 13 22 1 pmod w=100u l=10u
m21 22 13 23 1 pmod w=100u l=10u
m22 23 12 24 1 pmod w=100u l=10u
m23 24 11 1 1 pmod w=100u l=10u
m24 22 15 1 1 pmod w=100u l=10u
xc 15 26 1 inverter
xs 21 27 1 inverter
.tran 0.01ms 200ms
.control
run
plot V(11) V(12) V(13)
plot V(26) V(27)
.endc 
.end
