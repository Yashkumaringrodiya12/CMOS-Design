** DC Analysis
Vin 1 0 5.0
R1 1 2 0.5k
L1 2 3 100
C1 3 0 1u
.dc Vin 0.0 5.0 0.1
.control
run 
plot V(1) V(2)
.endc
.end