** Transient Analysis
Vin 1 0 pulse(0 5 0ns 0ns 0ns 100ms 200ms)
R1 1 2 8k
R2 2 0 2k
.tran 0.2ms 2000ms
.control
run 
plot V(1) V(2) 
.endc
.end
