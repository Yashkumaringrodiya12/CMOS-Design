** DC Analysis
Vin 1 0 5.0
R1 1 2 8k
R2 2 0 2k
.dc Vin 0.0 5.0 0.1
.control
run 
plot V(1) V(2)
.endc
.end