** DC Analysis
Vin 1 0 dc 0 ac 5
R1 1 2 8k
R2 2 0 16uF
.dc Vin 0.0 5.0 0.1
.control
run 
plot V(1) V(2)
.endc
.end